// 此文件描述的是指令集 irom 的设计
module irom(
    input clk,
    input [4:0]a,
    output reg [31:0]spo
);
    reg [31:0] strs [31:0]; // 32 λ��32��ָ��
    integer i_reg = 0;
    initial begin
        for(i_reg = 0; i_reg < 32; i_reg = i_reg + 1) begin
            strs[i_reg] = 32'h00000000;
        end
        strs[0] = 32'b00000000010000110010000000100000; // main: add $4, $2, $3
        strs[1] = 32'b10011100010001000000000000000100; //lw $4,4($2)
        strs[2] = 32'b10101100010001010000000000001000; //sw $5,8($2)
        strs[3] = 32'b00000000100000110001000000100010; // sub $2, $4, $3
        strs[4] = 32'b00000000100000110001000000100101;  //or $2,$4,$3
        strs[5] = 32'b00000000100000110001000000100100; // and $2, $4, $3
        strs[6] = 32'b00000000100000110001000000101010; //slt $2, $4, $3
        strs[7] = 32'b00001100000000000000000000000101; // jal addf
        strs[8] = 32'b00010000011000110000000000000001; //beq $3, $3, equ
        strs[9] = 32'b10011100011000100000000000000000; //lw $4,4($2)
        strs[10] = 32'b00010000100000110000000000000001; //equ : beq $3, $4, exit
        strs[11] = 32'b10101100011000100000000000000000; //sw $2,0($3)
        strs[12] = 32'b00001000000000000000000000000000; //exit : j main
        strs[13] = 32'b00000000101001010010100000100000; // addf: add $5, $5, $5
        strs[14] = 32'b00100000000000000000000000000000; //jr
    end
    always @(posedge clk) begin spo = strs[a]; end
endmodule

